// Copyright(C) 2021 Erdet Nasufi. All rights reserved.

module vsp
